--
-- VHDL Package Header work.util
--
-- Created:
--          by - bmarc.UNKNOWN (LAPTOP-TS0CSSEU)
--          at - 08:40:39 10/ 1/2020
--
-- using Mentor Graphics HDL Designer(TM) 2020.3 Built on 12 Jul 2020 at 11:01:26
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE pkg_util IS
END pkg_util;

PACKAGE BODY pkg_util IS
    
END PACKAGE BODY;